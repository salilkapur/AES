../AES.srcs/sources_1/new/gcm_aes.sv