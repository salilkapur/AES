../AES.srcs/sources_1/new/clk_gen.sv