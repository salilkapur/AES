../AES.srcs/sources_1/new/aes_encrypt.sv