../AES.srcs/sources_1/new/aes_encrypt_stage.sv