../AES.srcs/sim_1/imports/new/testbench.sv