../AES.srcs/sources_1/new/aes.sv